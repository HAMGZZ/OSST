-- THIS IS THE FIRST FILE?
