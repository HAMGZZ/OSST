-- PS/2 Driver PS/2 to ASCII