-- Main Top file
